** sch_path: /home/juandsr/PROJECTS/DAY1/xschem/INV_2_TB.sch
**.subckt INV_2_TB Vin Vout
*.opin Vin
*.opin Vout
x1 net1 Vin net2 GND INV_2
Vin Vin GND pulse(0 1.8 1ns 1ns 1ns 4ns 10ns)
.save i(vin)
V2 net1 GND 1.8
.save i(v2)
x2 net1 net2 net3 GND INV_16
x3 net1 net3 net4 GND INV_2
x4 net1 net4 net5 GND INV_16
x5 net1 net5 net6 GND INV_2
x6 net1 net6 Vout GND INV_16
**** begin user architecture code

** opencircuitdesign pdks install
.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt



.tran 0.0001n 50n
.save all

**** end user architecture code
**.ends

* expanding   symbol:  INV_2.sym # of pins=4
** sym_path: /home/juandsr/PROJECTS/DAY1/xschem/INV_2.sym
** sch_path: /home/juandsr/PROJECTS/DAY1/xschem/INV_2.sch
.subckt INV_2 VDD IN OUT VSS
*.ipin IN
*.opin OUT
*.iopin VDD
*.iopin VSS
XM1 OUT IN VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 OUT IN VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1.3 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  INV_16.sym # of pins=4
** sym_path: /home/juandsr/PROJECTS/DAY1/xschem/INV_16.sym
** sch_path: /home/juandsr/PROJECTS/DAY1/xschem/INV_16.sch
.subckt INV_16 VDD IN OUT VSS
*.ipin IN
*.opin OUT
*.iopin VDD
*.iopin VSS
XM1 OUT IN VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=16 nf=16 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 OUT IN VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=10.4 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
